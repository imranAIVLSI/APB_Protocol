module hw_top;


endmodule; hw_top